netcdf wind {
dimensions:
	bound = 2 ;
	lon = 10 ;
	lat = 10 ;
variables:
double lon(lon) ;
	lon:bounds = "lon_bnds" ;
	lon:units = "degree_east" ;
	lon:standard_name = "longitude" ;
double lon_bnds(lon, bound) ;
double lat(lat) ;
	lat:bounds = "lat_bnds" ;
	lat:units = "degree_north" ;
	lat:standard_name = "latitude" ;
double lat_bnds(lat, bound) ;
float wind_x-velocity(lat, lon) ;
	wind_x-velocity:coordinates = "lon lat" ;
	wind_x-velocity:units = "m s-1" ;
	wind_x-velocity:missing_value = -1.0E30 ;

// global attributes:
	:history = "Created Tue Apr 24 18:14:35 2018 by /Users/lemmen/devel/MOSSCO/code/scripts/create_gridspec.py" ;
	:creator = "Carsten Lemmen <carsten.lemmen@hzg.de>" ;
	:license = "Creative Commons share-alike (CCSA)" ;
	:copyright = "Helmholtz-Zentrum Geesthacht" ;
	:Conventions = "CF-1.6" ;

data:

 lon = 7.825, 7.875, 7.925, 7.975, 8.025, 8.075, 8.125, 8.175, 8.225, 8.275 ;

 lon_bnds =
  7.8, 7.85,
  7.85, 7.9,
  7.9, 7.95,
  7.95, 8,
  8, 8.05,
  8.05, 8.1,
  8.1, 8.15,
  8.15, 8.2,
  8.2, 8.25,
  8.25, 8.3 ;

 lat = 54.4915, 54.4945, 54.4975, 54.5005, 54.5035, 54.5065, 54.5095,
    54.5125, 54.5155, 54.5185 ;

 lat_bnds =
  54.49, 54.493,
  54.493, 54.496,
  54.496, 54.499,
  54.499, 54.502,
  54.502, 54.505,
  54.505, 54.508,
  54.508, 54.511,
  54.511, 54.514,
  54.514, 54.517,
  54.517, 54.52 ;

 wind_x-velocity =
  0.7975118, 0.7976561, 0.7978011, 0.7979471, 0.798094, 0.7982417, 0.7983903,
    0.7985398, 0.7986901, 0.7988413,
  0.7975719, 0.7977161, 0.7978612, 0.7980072, 0.798154, 0.7983017, 0.7984503,
    0.7985997, 0.79875, 0.7989012,
  0.797632, 0.7977762, 0.7979212, 0.7980672, 0.798214, 0.7983617, 0.7985103,
    0.7986597, 0.7988099, 0.7989611,
  0.7976921, 0.7978362, 0.7979813, 0.7981272, 0.798274, 0.7984217, 0.7985702,
    0.7987196, 0.7988699, 0.799021,
  0.7977521, 0.7978963, 0.7980413, 0.7981872, 0.798334, 0.7984816, 0.7986302,
    0.7987795, 0.7989298, 0.7990809,
  0.7978122, 0.7979563, 0.7981013, 0.7982472, 0.798394, 0.7985416, 0.7986901,
    0.7988394, 0.7989897, 0.7991408,
  0.7978722, 0.7980164, 0.7981613, 0.7983072, 0.798454, 0.7986016, 0.79875,
    0.7988994, 0.7990496, 0.7992007,
  0.7979323, 0.7980764, 0.7982213, 0.7983672, 0.7985139, 0.7986615, 0.79881,
    0.7989593, 0.7991095, 0.7992606,
  0.7979923, 0.7981364, 0.7982814, 0.7984272, 0.7985739, 0.7987215,
    0.7988699, 0.7990192, 0.7991694, 0.7993205,
  0.7980524, 0.7981964, 0.7983414, 0.7984872, 0.7986339, 0.7987815,
    0.7989299, 0.7990791, 0.7992293, 0.7993803 ;
}
