netcdf particle_scrip {
dimensions:
	grid_size = 138 ;
	grid_corners = 4 ;
	grid_rank = 2 ;
variables:
	int grid_dims(grid_rank) ;
		grid_dims:units = "unitless" ;
	int grid_imask(grid_size) ;
		grid_imask:units = "unitless" ;
	double grid_center_lat(grid_size) ;
		grid_center_lat:units = "degrees" ;
	double grid_center_lon(grid_size) ;
		grid_center_lon:units = "degrees" ;
	double grid_corner_lat(grid_size, grid_corners) ;
		grid_corner_lat:units = "degrees" ;
	double grid_corner_lon(grid_size, grid_corners) ;
		grid_corner_lon:units = "degrees" ;

// global attributes:
		:history = "Created Tue Dec 19 18:25:04 2017 by /Users/lemmen/devel/MOSSCO/code/scripts/bdy2scrip.py" ;
		:creator = "Carsten Lemmen <carsten.lemmen@hzg.de>" ;
		:license = "Creative Commons Attribution Share-alike (CC-BY-SA)" ;
		:copyright = "Helmholtz-Zentrum Geesthacht" ;
		:Conventions = "SCRIP" ;
data:

 grid_dims = 138, 4 ;

 grid_imask = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 grid_center_lat = 51.258861541748, 51.2768859863281, 51.2949371337891, 
    51.3130187988281, 51.3311500549316, 51.3493347167969, 51.3675918579102, 
    51.3859252929688, 51.4043502807617, 51.4228744506836, 51.4415092468262, 
    51.4602661132812, 51.4791564941406, 51.4981842041016, 51.5173645019531, 
    51.5367050170898, 51.5562133789062, 51.5758972167969, 51.5957717895508, 
    51.615837097168, 51.6361045837402, 51.6565818786621, 51.6772766113281, 
    51.6981964111328, 51.719352722168, 51.7407417297363, 51.7623748779297, 
    51.7842636108398, 51.8064117431641, 51.8288192749023, 51.8514976501465, 
    51.8744506835938, 51.8976821899414, 51.9211959838867, 51.9450035095215, 
    51.9691009521484, 51.9934997558594, 52.0181999206543, 52.0432052612305, 
    52.0685195922852, 54.1537780761719, 54.2037544250488, 54.2516174316406, 
    54.2983207702637, 54.3443603515625, 54.3899917602539, 54.4354019165039, 
    54.4807434082031, 54.5261726379395, 54.5718841552734, 54.6182174682617, 
    54.6654586791992, 54.7067260742188, 54.745189666748, 54.7818756103516, 
    54.8175430297852, 54.8525543212891, 54.8871078491211, 54.9213523864746, 
    54.9554214477539, 54.9894561767578, 55.0237083435059, 55.0582160949707, 
    55.085823059082, 55.1105575561523, 55.1334915161133, 55.1554107666016, 
    55.1766204833984, 55.1972808837891, 55.2174987792969, 55.2373199462891, 
    55.2568130493164, 55.2760162353516, 55.2949600219727, 55.3136978149414, 
    55.3322677612305, 55.350772857666, 55.3668746948242, 55.3805885314941, 
    55.3931617736816, 55.4051132202148, 55.4166488647461, 55.427848815918, 
    55.4387741088867, 55.4494552612305, 55.4599075317383, 55.4701499938965, 
    55.4802017211914, 55.4900665283203, 55.4997634887695, 55.5093002319336, 
    55.5186767578125, 55.5279083251953, 55.5370025634766, 55.5447654724121, 
    55.5508499145508, 55.5562438964844, 55.5612640380859, 55.5660514831543, 
    55.5706481933594, 55.5750923156738, 55.5793914794922, 55.5835647583008, 
    55.5876159667969, 55.591552734375, 55.5953750610352, 55.5990905761719, 
    55.6027069091797, 55.6062240600586, 55.6096458435059, 55.6129722595215, 
    55.6162071228027, 55.6193542480469, 55.6224098205566, 55.6253814697266, 
    55.6282577514648, 55.631046295166, 55.6337356567383, 55.6362991333008, 
    55.6380081176758, 55.6383323669434, 55.6382637023926, 55.6379852294922, 
    55.6376037597656, 55.6371574401855, 55.6366653442383, 55.6361465454102, 
    55.6355972290039, 55.6350250244141, 55.6344337463379, 55.6338272094727, 
    55.6331939697266, 55.6325531005859, 55.631893157959, 55.6312141418457, 
    55.6305160522461, 55.6297988891602, 55.6290512084961 ;

 grid_center_lon = 2.90595769882202, 2.87709975242615, 2.84820771217346, 
    2.81925916671753, 2.79023313522339, 2.76110816001892, 2.73186469078064, 
    2.70248293876648, 2.67294406890869, 2.64322900772095, 2.61332011222839, 
    2.5831995010376, 2.55284976959229, 2.52225399017334, 2.4913957118988, 
    2.46025848388672, 2.42882704734802, 2.39708566665649, 2.36501884460449, 
    2.33261251449585, 2.29985189437866, 2.26672315597534, 2.23321223258972, 
    2.19930624961853, 2.16499185562134, 2.13025665283203, 2.09508848190308, 
    2.05947470664978, 2.02340412139893, 1.98686504364014, 1.94984686374664, 
    1.91233849525452, 1.87432956695557, 1.83581006526947, 1.79676997661591, 
    1.75719976425171, 1.71709012985229, 1.67643189430237, 1.63521647453308, 
    1.59343528747559, -0.152019649744034, -0.0541966110467911, 
    0.0430246032774448, 0.139455139636993, 0.235447555780411, 
    0.331331849098206, 0.427405834197998, 0.523974418640137, 
    0.621402621269226, 0.720214128494263, 0.821390509605408, 
    0.930269718170166, 1.04332256317139, 1.15494918823242, 1.26473808288574, 
    1.37312686443329, 1.48061811923981, 1.58762717247009, 1.69454169273376, 
    1.80179357528687, 1.90997087955475, 2.02013826370239, 2.13759207725525, 
    2.25755548477173, 2.37429237365723, 2.48775386810303, 2.59858989715576, 
    2.7073802947998, 2.81452465057373, 2.92031621932983, 3.02499198913574, 
    3.12875843048096, 3.23181676864624, 3.33438539505005, 3.43673801422119, 
    3.53929853439331, 3.64307117462158, 3.7502326965332, 3.85452580451965, 
    3.95636510848999, 4.05604314804077, 4.15395402908325, 4.25036239624023, 
    4.3454532623291, 4.43936538696289, 4.53221321105957, 4.62409114837646, 
    4.71508979797363, 4.80529499053955, 4.89480113983154, 4.98371601104736, 
    5.07218551635742, 5.16044044494629, 5.24899864196777, 5.33927536010742, 
    5.42728996276855, 5.51325654983521, 5.59736061096191, 5.67987012863159, 
    5.76096105575562, 5.84074878692627, 5.91931629180908, 5.99672508239746, 
    6.07302188873291, 6.14824867248535, 6.22243642807007, 6.29561614990234, 
    6.36781311035156, 6.43905258178711, 6.50936031341553, 6.57876110076904, 
    6.64728212356567, 6.7149543762207, 6.78181409835815, 6.84790754318237, 
    6.91329717636108, 6.97807264328003, 7.04238367080688, 7.10655498504639, 
    7.17170333862305, 7.2346658706665, 7.29568386077881, 7.35493946075439, 
    7.4126443862915, 7.46895360946655, 7.52397632598877, 7.57779550552368, 
    7.6304783821106, 7.6820821762085, 7.7326602935791, 7.78226089477539, 
    7.83093309402466, 7.87872409820557, 7.92568445205688, 7.9718656539917, 
    8.01732540130615, 8.0621280670166, 8.10635375976562 ;

 grid_corner_lat =
  51.229923248291, 51.2698249816895, 51.2877998352051, 51.2479782104492,
  51.2479782104492, 51.2877998352051, 51.3057975769043, 51.2660484313965,
  51.2660484313965, 51.3057975769043, 51.3238296508789, 51.2841377258301,
  51.2841377258301, 51.3238296508789, 51.3419036865234, 51.3022689819336,
  51.3022689819336, 51.3419036865234, 51.3600311279297, 51.320442199707,
  51.320442199707, 51.3600311279297, 51.3782272338867, 51.338680267334,
  51.338680267334, 51.3782272338867, 51.3964996337891, 51.3569869995117,
  51.3569869995117, 51.3964996337891, 51.4148635864258, 51.375373840332,
  51.375373840332, 51.4148635864258, 51.4333229064941, 51.393856048584,
  51.393856048584, 51.4333229064941, 51.4518890380859, 51.4124412536621,
  51.4124412536621, 51.4518890380859, 51.4705772399902, 51.4311408996582,
  51.4311408996582, 51.4705772399902, 51.4893913269043, 51.4499664306641,
  51.4499664306641, 51.4893913269043, 51.5083465576172, 51.468921661377,
  51.468921661377, 51.5083465576172, 51.5274467468262, 51.4880218505859,
  51.4880218505859, 51.5274467468262, 51.5467071533203, 51.5072784423828,
  51.5072784423828, 51.5467071533203, 51.5661315917969, 51.5266914367676,
  51.5266914367676, 51.5661315917969, 51.5857353210449, 51.5462799072266,
  51.5462799072266, 51.5857353210449, 51.6055183410645, 51.566047668457,
  51.566047668457, 51.6055183410645, 51.6254959106445, 51.5860023498535,
  51.5860023498535, 51.6254959106445, 51.6456718444824, 51.6061515808105,
  51.6061515808105, 51.6456718444824, 51.6660575866699, 51.6265068054199,
  51.6265068054199, 51.6660575866699, 51.6866569519043, 51.6470718383789,
  51.6470718383789, 51.6866569519043, 51.7074813842773, 51.6678581237793,
  51.6678581237793, 51.7074813842773, 51.7285385131836, 51.6888732910156,
  51.6888732910156, 51.7285385131836, 51.749828338623, 51.7101173400879,
  51.7101173400879, 51.749828338623, 51.7713661193848, 51.7316017150879,
  51.7316017150879, 51.7713661193848, 51.7931518554688, 51.7533340454102,
  51.7533340454102, 51.7931518554688, 51.8151931762695, 51.775318145752,
  51.775318145752, 51.8151931762695, 51.8375015258789, 51.7975616455078,
  51.7975616455078, 51.8375015258789, 51.8600769042969, 51.8200721740723,
  51.8200721740723, 51.8600769042969, 51.8829231262207, 51.842845916748,
  51.842845916748, 51.8829231262207, 51.9060516357422, 51.8658981323242,
  51.8658981323242, 51.9060516357422, 51.9294662475586, 51.8892288208008,
  51.8892288208008, 51.9294662475586, 51.9531669616699, 51.9128456115723,
  51.9128456115723, 51.9531669616699, 51.9771614074707, 51.9367523193359,
  51.9367523193359, 51.9771614074707, 52.0014533996582, 51.9609527587891,
  51.9609527587891, 52.0014533996582, 52.026050567627, 51.9854469299316,
  51.9854469299316, 52.026050567627, 52.050952911377, 52.0102462768555,
  52.0102462768555, 52.050952911377, 52.0761642456055, 52.0353469848633,
  52.0353469848633, 52.0761642456055, 52.1016883850098, 52.0607604980469,
  54.1029815673828, 54.1549263000488, 54.1506385803223, 0,
  54.1549263000488, 54.2038841247559, 54.2045783996582, 0,
  54.2038841247559, 54.2512054443359, 54.2525825500488, 0,
  54.2512054443359, 54.2975921630859, 54.2993469238281, 0,
  54.2975921630859, 54.343391418457, 54.3454360961914, 0,
  54.343391418457, 54.3888168334961, 54.3911247253418, 0,
  54.3888168334961, 54.4340209960938, 54.4365882873535, 0,
  54.4340209960938, 54.4791259765625, 54.4819869995117, 0,
  54.4791259765625, 54.5242500305176, 54.5274696350098, 0,
  54.5242500305176, 54.5694770812988, 54.5732192993164, 0,
  54.5694770812988, 54.6147384643555, 54.6195220947266, 0,
  54.6147384643555, 54.6587791442871, 54.6669616699219, 0,
  54.6587791442871, 54.6991767883301, 54.7161827087402, 0,
  54.6991767883301, 54.7369537353516, 54.7546730041504, 0,
  54.7369537353516, 54.773323059082, 54.791202545166, 0,
  54.773323059082, 54.8087882995605, 54.8267936706543, 0,
  54.8087882995605, 54.843620300293, 54.8617668151855, 0,
  54.843620300293, 54.8779754638672, 54.8963241577148, 0,
  54.8779754638672, 54.9119758605957, 54.9305992126465, 0,
  54.9119758605957, 54.9456939697266, 54.964729309082, 0,
  54.9456939697266, 54.9791717529297, 54.9988632202148, 0,
  54.9791717529297, 55.0122108459473, 55.0332221984863, 0,
  55.0122108459473, 55.0434303283691, 55.068244934082, 0,
  55.0434303283691, 55.0705146789551, 55.1042213439941, 0,
  55.0705146789551, 55.0948295593262, 55.1282119750977, 0,
  55.0948295593262, 55.1177139282227, 55.1506004333496, 0,
  55.1177139282227, 55.1396713256836, 55.1721534729004, 0,
  55.1396713256836, 55.1609382629395, 55.1931037902832, 0,
  55.1609382629395, 55.1816520690918, 55.2135696411133, 0,
  55.1816520690918, 55.2018928527832, 55.2336273193359, 0,
  55.2018928527832, 55.2217254638672, 55.2533416748047, 0,
  55.2217254638672, 55.2411994934082, 55.2727508544922, 0,
  55.2411994934082, 55.2603378295898, 55.2919006347656, 0,
  55.2603378295898, 55.2791709899902, 55.3108291625977, 0,
  55.2791709899902, 55.2976875305176, 55.3295822143555, 0,
  55.2976875305176, 55.3158187866211, 55.3482208251953, 0,
  55.3158187866211, 55.3331642150879, 55.3668441772461, 0,
  55.3331642150879, 55.348560333252, 55.3857269287109, 0,
  55.348560333252, 55.3621101379395, 55.4005851745605, 0,
  55.3621101379395, 55.3747406005859, 55.4126167297363, 0,
  55.3747406005859, 55.3868103027344, 55.4242134094238, 0,
  55.3868103027344, 55.3984603881836, 55.4354858398438, 0,
  55.3984603881836, 55.4097747802734, 55.4464836120605, 0,
  55.4097747802734, 55.4207954406738, 55.4572372436523, 0,
  55.4207954406738, 55.4315490722656, 55.4677772521973, 0,
  55.4315490722656, 55.4420623779297, 55.4781112670898, 0,
  55.4420623779297, 55.4523506164551, 55.4882621765137, 0,
  55.4523506164551, 55.4624252319336, 55.4982376098633, 0,
  55.4624252319336, 55.4722938537598, 55.5080490112305, 0,
  55.4722938537598, 55.4819602966309, 55.5177116394043, 0,
  55.4819602966309, 55.4914207458496, 55.5272369384766, 0,
  55.4914207458496, 55.500659942627, 55.5366363525391, 0,
  55.500659942627, 55.5096168518066, 55.5459327697754, 0,
  55.5096168518066, 55.5180511474609, 55.5551567077637, 0,
  55.5180511474609, 55.5253143310547, 55.5643882751465, 0,
  55.5253143310547, 55.5313873291016, 55.5714797973633, 0,
  55.5313873291016, 55.5368728637695, 55.5763893127441, 0,
  55.5368728637695, 55.5420227050781, 55.5811042785645, 0,
  55.5420227050781, 55.5469284057617, 55.5856590270996, 0,
  55.5469284057617, 55.5516395568848, 55.5900802612305, 0,
  55.5516395568848, 55.5561828613281, 55.5943717956543, 0,
  55.5561828613281, 55.5605697631836, 55.5985450744629, 0,
  55.5605697631836, 55.5648193359375, 55.6026039123535, 0,
  55.5648193359375, 55.5689353942871, 55.606559753418, 0,
  55.5689353942871, 55.572925567627, 55.6104125976562, 0,
  55.572925567627, 55.5767974853516, 55.6141662597656, 0,
  55.5767974853516, 55.5805511474609, 55.6178207397461, 0,
  55.5805511474609, 55.5841941833496, 55.6213874816895, 0,
  55.5841941833496, 55.5877304077148, 55.6248626708984, 0,
  55.5877304077148, 55.5911560058594, 55.6282539367676, 0,
  55.5911560058594, 55.5944786071777, 55.6315612792969, 0,
  55.5944786071777, 55.5976982116699, 55.6347885131836, 0,
  55.5976982116699, 55.6008071899414, 55.6379356384277, 0,
  55.6008071899414, 55.6038131713867, 55.6410102844238, 0,
  55.6038131713867, 55.6067008972168, 55.6440124511719, 0,
  55.6067008972168, 55.6094627380371, 55.6469459533691, 0,
  55.6094627380371, 55.6120719909668, 55.6498184204102, 0,
  55.6120719909668, 55.6144638061523, 55.6526298522949, 0,
  55.6144638061523, 55.6164703369141, 55.6553955078125, 0,
  55.6164703369141, 55.617733001709, 55.6581344604492, 0,
  55.617733001709, 55.6182098388672, 55.6595420837402, 0,
  55.6182098388672, 55.6182746887207, 55.6589317321777, 0,
  55.6182746887207, 55.6181411743164, 55.658317565918, 0,
  55.6181411743164, 55.6178970336914, 55.6576957702637, 0,
  55.6178970336914, 55.6175689697266, 55.6570625305176, 0,
  55.6175689697266, 55.6171875, 55.6564178466797, 0,
  55.6171875, 55.6167602539062, 55.6557655334473, 0,
  55.6167602539062, 55.6162948608398, 55.655101776123, 0,
  55.6162948608398, 55.615795135498, 55.6544342041016, 0,
  55.615795135498, 55.6152648925781, 55.6537590026855, 0,
  55.6152648925781, 55.6147041320801, 55.6530723571777, 0,
  55.6147041320801, 55.6141166687012, 55.6523857116699, 0,
  55.6141166687012, 55.6135025024414, 55.6516876220703, 0,
  55.6135025024414, 55.6128578186035, 55.6509895324707, 0,
  55.6128578186035, 55.6121826171875, 55.6502838134766, 0,
  55.6121826171875, 55.6114654541016, 55.6495704650879, 0,
  55.6114654541016, 55.6106986999512, 55.648853302002, 0,
  55.6106986999512, 55.6098670959473, 55.6481323242188, 0 ;

 grid_corner_lon =
  2.88860034942627, 2.9521963596344, 2.92331480979919, 2.85978531837463,
  2.85978531837463, 2.92331480979919, 2.89441418647766, 2.83094382286072,
  2.83094382286072, 2.89441418647766, 2.86547160148621, 2.80205345153809,
  2.80205345153809, 2.86547160148621, 2.83646512031555, 2.77309250831604,
  2.77309250831604, 2.83646512031555, 2.80737376213074, 2.74403977394104,
  2.74403977394104, 2.80737376213074, 2.7781765460968, 2.71487545967102,
  2.71487545967102, 2.7781765460968, 2.74885392189026, 2.68557929992676,
  2.68557929992676, 2.74885392189026, 2.7193865776062, 2.6561324596405,
  2.6561324596405, 2.7193865776062, 2.6897554397583, 2.62651610374451,
  2.62651610374451, 2.6897554397583, 2.65994191169739, 2.59671187400818,
  2.59671187400818, 2.65994191169739, 2.62992835044861, 2.56670165061951,
  2.56670165061951, 2.62992835044861, 2.59969711303711, 2.53646850585938,
  2.53646850585938, 2.59969711303711, 2.5692310333252, 2.50599479675293,
  2.50599479675293, 2.5692310333252, 2.53851294517517, 2.47526431083679,
  2.47526431083679, 2.53851294517517, 2.50752711296082, 2.44426012039185,
  2.44426012039185, 2.50752711296082, 2.47625708580017, 2.41296672821045,
  2.41296672821045, 2.47625708580017, 2.4446873664856, 2.38136839866638,
  2.38136839866638, 2.4446873664856, 2.41280293464661, 2.349449634552,
  2.349449634552, 2.41280293464661, 2.38058829307556, 2.31719565391541,
  2.31719565391541, 2.38058829307556, 2.34802937507629, 2.28459191322327,
  2.28459191322327, 2.34802937507629, 2.31511187553406, 2.25162410736084,
  2.25162410736084, 2.31511187553406, 2.28182196617126, 2.21827840805054,
  2.21827840805054, 2.28182196617126, 2.24814605712891, 2.18454122543335,
  2.18454122543335, 2.24814605712891, 2.21407127380371, 2.15039944648743,
  2.15039944648743, 2.21407127380371, 2.17958426475525, 2.1158401966095,
  2.1158401966095, 2.17958426475525, 2.14467334747314, 2.08085107803345,
  2.08085107803345, 2.14467334747314, 2.10932564735413, 2.04541945457458,
  2.04541945457458, 2.10932564735413, 2.07352995872498, 2.00953364372253,
  2.00953364372253, 2.07352995872498, 2.03727436065674, 1.97318232059479,
  1.97318232059479, 2.03727436065674, 2.00054788589478, 1.93635404109955,
  1.93635404109955, 2.00054788589478, 1.96333968639374, 1.89903771877289,
  1.89903771877289, 1.96333968639374, 1.92563915252686, 1.86122298240662,
  1.86122298240662, 1.92563915252686, 1.88743615150452, 1.82289946079254,
  1.82289946079254, 1.88743615150452, 1.8487206697464, 1.78405690193176,
  1.78405690193176, 1.8487206697464, 1.80948305130005, 1.74468576908112,
  1.74468576908112, 1.80948305130005, 1.7697137594223, 1.70477640628815,
  1.70477640628815, 1.7697137594223, 1.72940385341644, 1.66431963443756,
  1.66431963443756, 1.72940385341644, 1.68854427337646, 1.62330651283264,
  1.62330651283264, 1.68854427337646, 1.64712655544281, 1.58172833919525,
  1.58172833919525, 1.64712655544281, 1.60514223575592, 1.53957664966583,
  -0.163516029715538, -0.0677515119314194, -0.246045336127281, 0,
  -0.0677515119314194, 0.0290014203637838, -0.140523254871368, 0,
  0.0290014203637838, 0.12521006166935, -0.0406417138874531, 0,
  0.12521006166935, 0.221017524600029, 0.0570477843284607, 0,
  0.221017524600029, 0.316704034805298, 0.153700232505798, 0,
  0.316704034805298, 0.412544369697571, 0.249877572059631, 0,
  0.412544369697571, 0.50882089138031, 0.345959663391113, 0,
  0.50882089138031, 0.605860352516174, 0.442267268896103, 0,
  0.605860352516174, 0.704098761081696, 0.539128005504608, 0,
  0.704098761081696, 0.804221510887146, 0.636944949626923, 0,
  0.804221510887146, 0.907523989677429, 0.736329555511475, 0,
  0.907523989677429, 1.01600539684296, 0.838559567928314, 0,
  1.01600539684296, 1.1270956993103, 0.953015506267548, 0,
  1.1270956993103, 1.23691523075104, 1.07063984870911, 0,
  1.23691523075104, 1.34534406661987, 1.18280279636383, 0,
  1.34534406661987, 1.45281326770782, 1.29256081581116, 0,
  1.45281326770782, 1.55971813201904, 1.4009096622467, 0,
  1.55971813201904, 1.66642427444458, 1.50842297077179, 0,
  1.66642427444458, 1.77331781387329, 1.61553609371185, 0,
  1.77331781387329, 1.88087713718414, 1.72265923023224, 0,
  1.88087713718414, 1.98981118202209, 1.83026945590973, 0,
  1.98981118202209, 2.10137414932251, 1.93906462192535, 0,
  2.10137414932251, 2.21725988388062, 2.05046510696411, 0,
  2.21725988388062, 2.33428359031677, 2.17381000518799, 0,
  2.33428359031677, 2.44843339920044, 2.29785084724426, 0,
  2.44843339920044, 2.55986428260803, 2.4143009185791, 0,
  2.55986428260803, 2.66914367675781, 2.52707409858704, 0,
  2.66914367675781, 2.77668809890747, 2.63731527328491, 0,
  2.77668809890747, 2.88280534744263, 2.74561715126038, 0,
  2.88280534744263, 2.98773884773254, 2.85236096382141, 0,
  2.98773884773254, 3.0916965007782, 2.95782732963562, 0,
  3.0916965007782, 3.19487309455872, 3.06224489212036, 0,
  3.19487309455872, 3.2974681854248, 3.16582012176514, 0,
  3.2974681854248, 3.39971232414246, 3.26876068115234, 0,
  3.39971232414246, 3.50191044807434, 3.37130260467529, 0,
  3.50191044807434, 3.60453319549561, 3.47376346588135, 0,
  3.60453319549561, 3.70831370353699, 3.5766863822937, 0,
  3.70831370353699, 3.81277847290039, 3.68160891532898, 0,
  3.81277847290039, 3.91534018516541, 3.79215145111084, 0,
  3.91534018516541, 4.01566886901855, 3.89627313613892, 0,
  4.01566886901855, 4.11414337158203, 3.99739027023315, 0,
  4.11414337158203, 4.2110481262207, 4.09641742706299, 0,
  4.2110481262207, 4.30658388137817, 4.19376468658447, 0,
  4.30658388137817, 4.40089845657349, 4.28967618942261, 0,
  4.40089845657349, 4.49411106109619, 4.38432216644287, 0,
  4.49411106109619, 4.5863208770752, 4.47783279418945, 0,
  4.5863208770752, 4.67761754989624, 4.57031488418579, 0,
  4.67761754989624, 4.76808547973633, 4.66186141967773, 0,
  4.76808547973633, 4.85781240463257, 4.75256156921387, 0,
  4.85781240463257, 4.9468936920166, 4.84250450134277, 0,
  4.9468936920166, 5.03544664382935, 4.93178939819336, 0,
  5.03544664382935, 5.12362957000732, 5.02053833007812, 0,
  5.12362957000732, 5.2116847038269, 5.10892486572266, 0,
  5.2116847038269, 5.29997253417969, 5.19725179672241, 0,
  5.29997253417969, 5.38825559616089, 5.28631210327148, 0,
  5.38825559616089, 5.47494983673096, 5.37857818603516, 0,
  5.47494983673096, 5.55973100662231, 5.46632385253906, 0,
  5.55973100662231, 5.64285326004028, 5.55156326293945, 0,
  5.64285326004028, 5.72451066970825, 5.63499069213867, 0,
  5.72451066970825, 5.80483150482178, 5.7168869972229, 0,
  5.80483150482178, 5.88390636444092, 5.79741144180298, 0,
  5.88390636444092, 5.96180200576782, 5.87666654586792, 0,
  5.96180200576782, 6.03857040405273, 5.9547266960144, 0,
  6.03857040405273, 6.11425447463989, 6.03164768218994, 0,
  6.11425447463989, 6.18888854980469, 6.10747385025024, 0,
  6.18888854980469, 6.26250314712524, 6.18224239349365, 0,
  6.26250314712524, 6.33512544631958, 6.25598430633545, 0,
  6.33512544631958, 6.40678071975708, 6.32872867584229, 0,
  6.40678071975708, 6.47749328613281, 6.40050029754639, 0,
  6.47749328613281, 6.547287940979, 6.4713249206543, 0,
  6.547287940979, 6.61618900299072, 6.5412278175354, 0,
  6.61618900299072, 6.68422603607178, 6.61023473739624, 0,
  6.68422603607178, 6.75143003463745, 6.67837524414062, 0,
  6.75143003463745, 6.81784009933472, 6.74568271636963, 0,
  6.81784009933472, 6.88350582122803, 6.81219816207886, 0,
  6.88350582122803, 6.94849252700806, 6.87797498703003, 0,
  6.94849252700806, 7.01289176940918, 6.94308853149414, 0,
  7.01289176940918, 7.07683801651001, 7.007652759552, 0,
  7.07683801651001, 7.14048528671265, 7.07187557220459, 0,
  7.14048528671265, 7.20363187789917, 7.13627243041992, 0,
  7.20363187789917, 7.26535415649414, 7.20292091369629, 0,
  7.26535415649414, 7.3253173828125, 7.265700340271, 0,
  7.3253173828125, 7.3836784362793, 7.32601356506348, 0,
  7.3836784362793, 7.44059944152832, 7.38456201553345, 0,
  7.44059944152832, 7.49619674682617, 7.44161033630371, 0,
  7.49619674682617, 7.55055999755859, 7.49730777740479, 0,
  7.55055999755859, 7.603759765625, 7.55175542831421, 0,
  7.603759765625, 7.65585517883301, 7.60503101348877, 0,
  7.65585517883301, 7.70690107345581, 7.65719699859619, 0,
  7.70690107345581, 7.75694608688354, 7.70830917358398, 0,
  7.75694608688354, 7.80603837966919, 7.75841951370239, 0,
  7.80603837966919, 7.85422468185425, 7.80757617950439, 0,
  7.85422468185425, 7.9015531539917, 7.85582780838013, 0,
  7.9015531539917, 7.94807291030884, 7.90322399139404, 0,
  7.94807291030884, 7.99383640289307, 7.94981575012207, 0,
  7.99383640289307, 8.03890037536621, 7.99565839767456, 0,
  8.03890037536621, 8.08332920074463, 8.04081439971924, 0,
  8.08332920074463, 8.12719440460205, 8.08535671234131, 0 ;
}
