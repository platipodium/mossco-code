netcdf wind {
dimensions:
	bound = 2 ;
	lon = 8 ;
	lat = 10 ;
variables:
	double lon(lon) ;
		lon:bounds = "lon_bnds" ;
		lon:units = "degree_east" ;
		lon:standard_name = "longitude" ;
	double lon_bnds(lon, bound) ;
	double lat(lat) ;
		lat:bounds = "lat_bnds" ;
		lat:units = "degree_north" ;
		lat:standard_name = "latitude" ;
	double lat_bnds(lat, bound) ;
	float wind_x-velocity(lat, lon) ;
		wind_x-velocity:coordinates = "lon lat" ;
		wind_x-velocity:units = "m s-1" ;

// global attributes:
		:history = "Created Tue Apr 24 18:14:35 2018 by /Users/lemmen/devel/MOSSCO/code/scripts/create_gridspec.py" ;
		:creator = "Carsten Lemmen <carsten.lemmen@hzg.de>" ;
		:license = "Creative Commons share-alike (CCSA)" ;
		:copyright = "Helmholtz-Zentrum Geesthacht" ;
		:Conventions = "CF-1.6" ;
data:

 lon = -12.5, -7.5, -2.5, 2.5, 7.5, 12.5, 17.5, 22.5 ;

 lon_bnds =
  -15, -10,
  -10, -5,
  -5, 0,
  0, 5,
  5, 10,
  10, 15,
  15, 20,
  20, 25 ;

 lat = 41.25, 43.75, 46.25, 48.75, 51.25, 53.75, 56.25, 58.75, 61.25, 63.75 ;

 lat_bnds =
  40, 42.5,
  42.5, 45,
  45, 47.5,
  47.5, 50,
  50, 52.5,
  52.5, 55,
  55, 57.5,
  57.5, 60,
  60, 62.5,
  62.5, 65 ;

 wind_x-velocity =
 0.5361943, 0.510237, 0.4970792, 0.4970792, 0.510237, 0.5361943, 0.5741901,
	 0.6229734,
 0.5896725, 0.5648005, 0.5521666, 0.5521666, 0.5648005, 0.5896725,
	 0.6259475, 0.6722689,
 0.6435996, 0.6199903, 0.6079686, 0.6079686, 0.6199903, 0.6435996,
	 0.6778871, 0.7213906,
 0.6972392, 0.6750829, 0.6637686, 0.6637686, 0.6750829, 0.6972392,
	 0.7292542, 0.7695619,
 0.7497559, 0.7292542, 0.7187485, 0.7187485, 0.7292542, 0.7497559,
	 0.7791983, 0.8159146,
 0.800216, 0.7815793, 0.7719879, 0.7719879, 0.7815793, 0.800216, 0.8267736,
	 0.8594901,
 0.8475889, 0.8310335, 0.8224657, 0.8224657, 0.8310335, 0.8475889,
	 0.8709428, 0.8992453,
 0.8907545, 0.876499, 0.8690654, 0.8690654, 0.876499, 0.8907545, 0.9105842,
	 0.9340603,
 0.928513, 0.9167736, 0.9105842, 0.9105842, 0.9167736, 0.928513, 0.9445037,
	 0.9627524,
 0.959601, 0.9505863, 0.9457477, 0.9457477, 0.9505863, 0.959601, 0.9714512,
	 0.9840934 ;
}
